`default_nettype none
`timescale 1ns / 1ps

/**
 * This is a PicoBlaze program memory.
 */
module ProgramMemory (
		
		/** the clock signal **/
		input clk,
		
		/** the current instruction address **/
		input [9:0] address,
		
		/** the instruction **/
		output [17:0] instruction
		
	);
	
	RAMB16_S18 blockRam(
		.DI (16'h0000),
		.DIP (2'b00),
		.EN (1'b1),
		.WE (1'b0),
		.SSR (1'b0),
		.CLK (clk),
		.ADDR (address),
		.DO (instruction[15:0]),
		.DOP (instruction[17:16])
	/*synthesis
init_00 = "0000000000000000000000000000000000000000000000000000000000004000"
init_01 = "0000000000000000000000000000000000000000000000000000000000000000"
init_02 = "0000000000000000000000000000000000000000000000000000000000000000"
init_03 = "0000000000000000000000000000000000000000000000000000000000000000"
init_04 = "0000000000000000000000000000000000000000000000000000000000000000"
init_05 = "0000000000000000000000000000000000000000000000000000000000000000"
init_06 = "0000000000000000000000000000000000000000000000000000000000000000"
init_07 = "0000000000000000000000000000000000000000000000000000000000000000"
init_08 = "0000000000000000000000000000000000000000000000000000000000000000"
init_09 = "0000000000000000000000000000000000000000000000000000000000000000"
init_0A = "0000000000000000000000000000000000000000000000000000000000000000"
init_0B = "0000000000000000000000000000000000000000000000000000000000000000"
init_0C = "0000000000000000000000000000000000000000000000000000000000000000"
init_0D = "0000000000000000000000000000000000000000000000000000000000000000"
init_0E = "0000000000000000000000000000000000000000000000000000000000000000"
init_0F = "0000000000000000000000000000000000000000000000000000000000000000"
init_10 = "0000000000000000000000000000000000000000000000000000000000000000"
init_11 = "0000000000000000000000000000000000000000000000000000000000000000"
init_12 = "0000000000000000000000000000000000000000000000000000000000000000"
init_13 = "0000000000000000000000000000000000000000000000000000000000000000"
init_14 = "0000000000000000000000000000000000000000000000000000000000000000"
init_15 = "0000000000000000000000000000000000000000000000000000000000000000"
init_16 = "0000000000000000000000000000000000000000000000000000000000000000"
init_17 = "0000000000000000000000000000000000000000000000000000000000000000"
init_18 = "0000000000000000000000000000000000000000000000000000000000000000"
init_19 = "0000000000000000000000000000000000000000000000000000000000000000"
init_1A = "0000000000000000000000000000000000000000000000000000000000000000"
init_1B = "0000000000000000000000000000000000000000000000000000000000000000"
init_1C = "0000000000000000000000000000000000000000000000000000000000000000"
init_1D = "0000000000000000000000000000000000000000000000000000000000000000"
init_1E = "0000000000000000000000000000000000000000000000000000000000000000"
init_1F = "0000000000000000000000000000000000000000000000000000000000000000"
init_20 = "0000000000000000000000000000000000000000000000000000000000000000"
init_21 = "0000000000000000000000000000000000000000000000000000000000000000"
init_22 = "0000000000000000000000000000000000000000000000000000000000000000"
init_23 = "0000000000000000000000000000000000000000000000000000000000000000"
init_24 = "0000000000000000000000000000000000000000000000000000000000000000"
init_25 = "0000000000000000000000000000000000000000000000000000000000000000"
init_26 = "0000000000000000000000000000000000000000000000000000000000000000"
init_27 = "0000000000000000000000000000000000000000000000000000000000000000"
init_28 = "0000000000000000000000000000000000000000000000000000000000000000"
init_29 = "0000000000000000000000000000000000000000000000000000000000000000"
init_2A = "0000000000000000000000000000000000000000000000000000000000000000"
init_2B = "0000000000000000000000000000000000000000000000000000000000000000"
init_2C = "0000000000000000000000000000000000000000000000000000000000000000"
init_2D = "0000000000000000000000000000000000000000000000000000000000000000"
init_2E = "0000000000000000000000000000000000000000000000000000000000000000"
init_2F = "0000000000000000000000000000000000000000000000000000000000000000"
init_30 = "0000000000000000000000000000000000000000000000000000000000000000"
init_31 = "0000000000000000000000000000000000000000000000000000000000000000"
init_32 = "0000000000000000000000000000000000000000000000000000000000000000"
init_33 = "0000000000000000000000000000000000000000000000000000000000000000"
init_34 = "0000000000000000000000000000000000000000000000000000000000000000"
init_35 = "0000000000000000000000000000000000000000000000000000000000000000"
init_36 = "0000000000000000000000000000000000000000000000000000000000000000"
init_37 = "0000000000000000000000000000000000000000000000000000000000000000"
init_38 = "0000000000000000000000000000000000000000000000000000000000000000"
init_39 = "0000000000000000000000000000000000000000000000000000000000000000"
init_3A = "0000000000000000000000000000000000000000000000000000000000000000"
init_3B = "0000000000000000000000000000000000000000000000000000000000000000"
init_3C = "0000000000000000000000000000000000000000000000000000000000000000"
init_3D = "0000000000000000000000000000000000000000000000000000000000000000"
init_3E = "0000000000000000000000000000000000000000000000000000000000000000"
init_3F = "0000000000000000000000000000000000000000000000000000000000000000"
initp_00 = "0000000000000000000000000000000000000000000000000000000000000003"
initp_01 = "0000000000000000000000000000000000000000000000000000000000000000"
initp_02 = "0000000000000000000000000000000000000000000000000000000000000000"
initp_03 = "0000000000000000000000000000000000000000000000000000000000000000"
initp_04 = "0000000000000000000000000000000000000000000000000000000000000000"
initp_05 = "0000000000000000000000000000000000000000000000000000000000000000"
initp_06 = "0000000000000000000000000000000000000000000000000000000000000000"
initp_07 = "0000000000000000000000000000000000000000000000000000000000000000"
*/);

// synthesis translate_off
defparam blockRam.INIT_00 = 256'h0000000000000000000000000000000000000000000000000000000000004000;
defparam blockRam.INIT_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_08 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_09 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_0A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_0B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_0C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_0D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_0E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_0F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_10 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_11 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_12 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_13 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_14 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_15 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_16 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_17 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_18 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_19 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_1A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_1B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_1C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_1D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_1E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_1F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_20 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_21 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_22 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_23 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_24 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_25 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_26 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_27 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_28 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_29 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_2A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_2B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_2C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_2D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_2E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_2F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_30 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_31 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_32 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_33 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_34 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_35 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_36 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_37 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_38 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_39 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_3A = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_3B = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_3C = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_3D = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_3E = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INIT_3F = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INITP_00 = 256'h0000000000000000000000000000000000000000000000000000000000000003;
defparam blockRam.INITP_01 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INITP_02 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INITP_03 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INITP_04 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INITP_05 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INITP_06 = 256'h0000000000000000000000000000000000000000000000000000000000000000;
defparam blockRam.INITP_07 = 256'h0000000000000000000000000000000000000000000000000000000000000000;

// synthesis translate_on
// synthesis attribute INIT_00 of blockRam is "0000000000000000000000000000000000000000000000000000000000004000"
// synthesis attribute INIT_01 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_02 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_03 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_04 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_05 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_06 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_07 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_08 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_09 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0A of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0B of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0C of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0D of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0E of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_0F of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_10 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_11 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_12 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_13 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_14 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_15 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_16 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_17 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_18 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_19 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1A of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1B of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1C of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1D of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1E of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_1F of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_20 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_21 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_22 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_23 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_24 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_25 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_26 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_27 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_28 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_29 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2A of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2B of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2C of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2D of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2E of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_2F of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_30 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_31 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_32 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_33 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_34 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_35 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_36 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_37 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_38 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_39 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3A of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3B of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3C of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3D of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3E of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INIT_3F of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INITP_00 of blockRam is "0000000000000000000000000000000000000000000000000000000000000003"
// synthesis attribute INITP_01 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INITP_02 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INITP_03 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INITP_04 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INITP_05 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INITP_06 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"
// synthesis attribute INITP_07 of blockRam is "0000000000000000000000000000000000000000000000000000000000000000"

endmodule

