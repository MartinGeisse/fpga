
module through(dataIn, ledOut);
	input dataIn;
	output ledOut;

	assign ledOut = dataIn;

endmodule
